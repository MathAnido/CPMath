module SL2(_input, output_);
	input [31:0] _input;		//Entrada do dado
	output reg [31:0] output_;	//Saida do dado
	always @ (*) begin
		output_ <= _input << 2;	//Atribuindo entrada deslocada em 2 bits na saida
	end	
endmodule
